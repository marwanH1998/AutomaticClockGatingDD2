

module test32bit
(
  D_IN,
  CLK,
  EN,
  D_OUT
);

  wire __clockgate_output_gclk_;
  wire [31:0] _00_;
  input CLK;
  input [31:0] D_IN;
  output [31:0] D_OUT;
  input EN;

  sky130_fd_sc_hd__dlclkp
  __clockgate_cell__
  (
    .GCLK(__clockgate_output_gclk_),
    .GATE(EN),
    .CLK(CLK)
  );


  sky130_fd_sc_hd__dfxtp_1
  _33_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[8]),
    .Q(D_OUT[8])
  );


  sky130_fd_sc_hd__dfxtp_1
  _34_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[13]),
    .Q(D_OUT[13])
  );


  sky130_fd_sc_hd__dfxtp_1
  _35_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[9]),
    .Q(D_OUT[9])
  );


  sky130_fd_sc_hd__dfxtp_1
  _36_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[6]),
    .Q(D_OUT[6])
  );


  sky130_fd_sc_hd__dfxtp_1
  _37_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[17]),
    .Q(D_OUT[17])
  );


  sky130_fd_sc_hd__dfxtp_1
  _38_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[26]),
    .Q(D_OUT[26])
  );


  sky130_fd_sc_hd__dfxtp_1
  _39_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[22]),
    .Q(D_OUT[22])
  );


  sky130_fd_sc_hd__dfxtp_1
  _40_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[27]),
    .Q(D_OUT[27])
  );


  sky130_fd_sc_hd__dfxtp_1
  _41_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[11]),
    .Q(D_OUT[11])
  );


  sky130_fd_sc_hd__dfxtp_1
  _42_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[10]),
    .Q(D_OUT[10])
  );


  sky130_fd_sc_hd__dfxtp_1
  _43_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[21]),
    .Q(D_OUT[21])
  );


  sky130_fd_sc_hd__dfxtp_1
  _44_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[16]),
    .Q(D_OUT[16])
  );


  sky130_fd_sc_hd__dfxtp_1
  _45_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[12]),
    .Q(D_OUT[12])
  );


  sky130_fd_sc_hd__dfxtp_1
  _46_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[25]),
    .Q(D_OUT[25])
  );


  sky130_fd_sc_hd__dfxtp_1
  _47_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[31]),
    .Q(D_OUT[31])
  );


  sky130_fd_sc_hd__dfxtp_1
  _48_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[24]),
    .Q(D_OUT[24])
  );


  sky130_fd_sc_hd__dfxtp_1
  _49_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[0]),
    .Q(D_OUT[0])
  );


  sky130_fd_sc_hd__dfxtp_1
  _50_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[3]),
    .Q(D_OUT[3])
  );


  sky130_fd_sc_hd__dfxtp_1
  _51_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[7]),
    .Q(D_OUT[7])
  );


  sky130_fd_sc_hd__dfxtp_1
  _52_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[4]),
    .Q(D_OUT[4])
  );


  sky130_fd_sc_hd__dfxtp_1
  _53_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[5]),
    .Q(D_OUT[5])
  );


  sky130_fd_sc_hd__dfxtp_1
  _54_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[2]),
    .Q(D_OUT[2])
  );


  sky130_fd_sc_hd__dfxtp_1
  _55_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[1]),
    .Q(D_OUT[1])
  );


  sky130_fd_sc_hd__dfxtp_1
  _56_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[23]),
    .Q(D_OUT[23])
  );


  sky130_fd_sc_hd__dfxtp_1
  _57_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[18]),
    .Q(D_OUT[18])
  );


  sky130_fd_sc_hd__dfxtp_1
  _58_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[15]),
    .Q(D_OUT[15])
  );


  sky130_fd_sc_hd__dfxtp_1
  _59_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[20]),
    .Q(D_OUT[20])
  );


  sky130_fd_sc_hd__dfxtp_1
  _60_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[19]),
    .Q(D_OUT[19])
  );


  sky130_fd_sc_hd__dfxtp_1
  _61_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[30]),
    .Q(D_OUT[30])
  );


  sky130_fd_sc_hd__dfxtp_1
  _62_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[28]),
    .Q(D_OUT[28])
  );


  sky130_fd_sc_hd__dfxtp_1
  _63_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[29]),
    .Q(D_OUT[29])
  );


  sky130_fd_sc_hd__dfxtp_1
  _64_
  (
    .CLK(__clockgate_output_gclk_),
    .D(D_IN[14]),
    .Q(D_OUT[14])
  );


endmodule

